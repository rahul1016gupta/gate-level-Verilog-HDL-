`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/30/2025 10:17:28 AM
// Design Name: 
// Module Name: ANDGATE_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ANDGATE_tb;
    reg A;
    reg B;
    wire Y;
AND_GATE dut(A,B,Y)
initial begin
A=1; B= 
    
    
endmodule
